module CLA_4bit(A, B, Cin, S, P, G, Ovfl);
input [3:0] A;
input [3:0] B;
output[3:0] S;
input Cin;
output P, G, Ovfl;

wire cout;
wire c1;
wire c2;
wire c3;
wire p0;
wire p1;
wire p2;
wire p3;
wire g0;
wire g1;
wire g2;
wire g3;

cla add_0(.A(A[0]), .B(B[0]), .C(Cin), .S(S[0]), .P(p0), .G(g0));
cla add_1(.A(A[1]), .B(B[1]), .C(c1), .S(S[1]), .P(p1), .G(g1));
cla add_2(.A(A[2]), .B(B[2]), .C(c2), .S(S[2]), .P(p2), .G(g2));
cla add_3(.A(A[3]), .B(B[3]), .C(c3), .S(S[3]), .P(p3), .G(g3));

assign c1 = g0 | (p0 &  Cin);
assign c2 = g1 | (g0 & p1) | (Cin & p0 & p1);
assign c3 = g2 | (g1 & p2) | (g0 & p1 & p2) | (Cin & p0 & p1 & p2);
assign cout = g3 | (g2 & p3) | (g1 & p2 & p3) | (g0 & p1 & p2 & p3) | (Cin & p0 & p1 & p2 & p3);

assign P = p0 & p1 & p2 & p3;
assign G = g3 | (g2 & p3) | (g1 & p2 & p3) | (g0 & p1 & p2 & p3);





endmodule
